library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity controller is
    port(
        instruction : in  std_logic_vector(15 downto 0);
        rst         : in  std_logic;
        pc_sel      : out std_logic;
        we_pc       : out std_logic;
        we_reg      : out std_logic;
        we_mem      : out std_logic;
        alu_sel_a   : out std_logic;
        alu_sel_b   : out std_logic_vector(1 downto 0);
        alu_opr     : out std_logic_vector(2 downto 0);
        wd_sel      : out std_logic
    );
end controller;

architecture Behavioral of controller is
    signal opcode : std_logic_vector(2 downto 0);
begin
    opcode <= instruction(15 downto 13);

    process(opcode, rst)
    begin
        if rst = '1' then
            pc_sel   <= '0';
            we_pc    <= '0';
            we_reg   <= '0';
            we_mem   <= '0';
            alu_sel_a <= '0';
            alu_sel_b <= "00";
            alu_opr  <= "000";
            wd_sel   <= '0';
        else
            case opcode is
                -- NEG: rA <- 2?s Complement (rB)
                when "000" =>
                    pc_sel   <= '0';
                    we_pc    <= '1';
                    we_reg   <= '1';
                    we_mem   <= '0';
                    alu_sel_a <= '1';
                    alu_sel_b <= "01";
                    alu_opr  <= "001";
                    wd_sel   <= '1';

                -- SBR: rB(Imm) <- ?1?
                when "001" =>
                    pc_sel   <= '0';
                    we_pc    <= '1';
                    we_reg   <= '1';
                    we_mem   <= '0';
                    alu_sel_a <= '0';
                    alu_sel_b <= "11";
                    alu_opr  <= "010";
                    wd_sel   <= '0';

                -- OR: rA <- [rB OR Z.F.(Imm)]
                when "010" =>
                    pc_sel   <= '0';
                    we_pc    <= '1';
                    we_reg   <= '1';
                    we_mem   <= '0';
                    alu_sel_a <= '1';
                    alu_sel_b <= "11";
                    alu_opr  <= "011";
                    wd_sel   <= '1';

                -- RJMP: PC <- 2*[PC + rA + S.E.(Imm)]
                when "011" =>
                    pc_sel   <= '1';
                    we_pc    <= '1';
                    we_reg   <= '0';
                    we_mem   <= '0';
                    alu_sel_a <= '1';
                    alu_sel_b <= "01";
                    alu_opr  <= "100";
                    wd_sel   <= '0';

                -- LUI: rA <- Imm * 128
                when "100" =>
                    pc_sel   <= '0';
                    we_pc    <= '1';
                    we_reg   <= '1';
                    we_mem   <= '0';
                    alu_sel_a <= '0';
                    alu_sel_b <= "11";
                    alu_opr  <= "101";
                    wd_sel   <= '1';

                -- LDI: rA <- Mem[2*Z.F.(Imm)]
                when "101" =>
                    pc_sel   <= '0';
                    we_pc    <= '1';
                    we_reg   <= '1';
                    we_mem   <= '0';
                    alu_sel_a <= '0';
                    alu_sel_b <= "11";
                    alu_opr  <= "110";
                    wd_sel   <= '0';

                -- STI: Mem[2*Z.F.(Imm)] <- rA
                when "110" =>
                    pc_sel   <= '0';
                    we_pc    <= '1';
                    we_reg   <= '0';
                    we_mem   <= '1';
                    alu_sel_a <= '1';
                    alu_sel_b <= "11";
                    alu_opr  <= "111";
                    wd_sel   <= '0';

                when others =>
                    pc_sel   <= '0';
                    we_pc    <= '0';
                    we_reg   <= '0';
                    we_mem   <= '0';
                    alu_sel_a <= '0';
                    alu_sel_b <= "00";
                    alu_opr  <= "000";
                    wd_sel   <= '0';
            end case;
        end if;
    end process;
end Behavioral;

